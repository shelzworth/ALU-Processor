LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY ssegmodified IS
PORT (
negative : IN STD_LOGIC;
bcd : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
leds, ledss: OUT STD_LOGIC_VECTOR(0 TO 6)
);
END ssegmodified;

ARCHITECTURE Behavior OF ssegmodified IS
BEGIN
PROCESS (bcd)
BEGIN
if negative = '1' then
ledss <= "1111110";
else
ledss <= "1111111";

END if;

CASE bcd IS   -- abcdefg
WHEN "0000" => leds <= "1101010";
WHEN "0001" => leds <= "1000100";
WHEN "0010" => leds <= "1101010";
WHEN "0011" => leds <= "1000100";
WHEN "0100" => leds <= "1101010";
WHEN "0101" => leds <= "1000100";
WHEN "0110" => leds <= "1101010";
WHEN "0111" => leds <= "1000100";
WHEN "1000" => leds <= "1101010";
WHEN "1001" => leds <= "1000100";
WHEN "1010" => leds <= "1101010";
WHEN "1011" => leds <= "1000100";
WHEN "1100" => leds <= "1101010";
WHEN "1101" => leds <= "1000100";
WHEN "1110" => leds <= "1101010";
WHEN "1111" => leds <= "1000100";
WHEN OTHERS => leds <= "-------";
END CASE;
END PROCESS;
END Behavior;
